module controlor(
    
);

endmodule // 控制器